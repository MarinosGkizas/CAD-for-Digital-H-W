module leds(x,s);
 input [3:0] x;
 output [9:0] s;

 assign s = (x == 4'd0 ) ? 10'b0000000001 :
 (x == 4'd1 ) ? 10'b0000000010 :
 (x == 4'd2 ) ? 10'b0000000100 : 
 (x == 4'd3 ) ? 10'b0000001000 :
 (x == 4'd4 ) ? 10'b0000010000 : 
 (x == 4'd5 ) ? 10'b0000100000 :
 (x == 4'd6 ) ? 10'b0001000000 : 
 (x == 4'd7 ) ? 10'b0010000000 :
 (x == 4'd8 ) ? 10'b0100000000 : 10'b1000000000 ;
 
 
endmodule